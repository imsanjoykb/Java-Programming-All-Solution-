* C:\Users\Sanjoy Kumar\Documents\JFETCdamplifier.sch

* Schematics Version 9.2
* Wed Jan 31 04:42:26 2018



** Analysis setup **
.DC LIN V_VDD 20 100 .01 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "JFETCdamplifier.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
