* C:\Users\Sanjoy Kumar\Documents\CurrentShuntfeedback.sch

* Schematics Version 9.2
* Wed Jan 31 04:26:22 2018



** Analysis setup **
.ac DEC 20 10 1Mhz
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "CurrentShuntfeedback.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
