* C:\Users\Sanjoy Kumar\Documents\Mosfetintegreted.sch

* Schematics Version 9.2
* Wed Jan 31 04:51:12 2018



** Analysis setup **
.DC LIN V_V1 10 100 .1 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Mosfetintegreted.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
